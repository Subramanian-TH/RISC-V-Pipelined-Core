module PC_Adder(
input [31:0] a, b,
output [31:0] r
    );
    
    assign r = a + b;
    
endmodule
